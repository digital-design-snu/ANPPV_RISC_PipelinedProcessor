`timescale 1ns / 1ps

 module MultiPortMem(
    input   [15:0]   addressInst,    // Address In :: Instruction Fetch address input :: PC
    input   [15:0]   addressOper,    // Address In :: Operand Fetch address input :: AS1
    input   [15:0]   addressWb,      // Address In :: WriteBack address input :: AS2
    input   [15:0]   dataWb,         // Data IN  :: From WriteBack Stage
    output  [15:0]   dataInst,       // Data OUT :: Instruction Fetch DataPath
    output  [15:0]   dataOper,       // Data OUT :: Operand Fetch Data Path
    input           writeEn,        // EN :: Write Enable From Write Back Stage
    input           clk             // Global Clock
    );
    reg  [15:0] blockMem[255:0];
    wire [15:0] addrPort2;
    // the code below avoids Write After Read Errors
    // Check Write Enable , if any read add  ==  write address then return vaalue in write bus to read bbus :? B)
    assign addrPort2 = (writeEn == 1'b1)? addressWb : addressOper ;
    assign dataInst = (writeEn&&(addrPort2 == addressInst))? dataWb : blockMem[addressInst]; 
    //assign dataOper = (writeEn&&(addressWb == addressOper))? dataWb : blockMem[addressOper];  // This Is useless now
    assign dataOper = blockMem[addrPort2] ;   
    
    always@(posedge clk) begin
        if(writeEn)
            blockMem[addrPort2] <= dataWb;
    end
 
    initial begin
    /*blockMem[0] = 8'h01; //CLR
    blockMem[1] = 8'h8;  //JCD<fl><od>
    blockMem[2] = 8'hc;  //JCD<fl><od>
    blockMem[3] = 8'h31;  //CCD<fl><od>
    blockMem[4] = 8'hd1;  //ORA<rn>
    blockMem[5] = 8'h79;  //POP<rn>
    blockMem[6] = 8'h2d;  //JCA<fl>
    blockMem[7] = 8'hc3;  //ANA<rn>
    blockMem[8] = 8'h4c;  //RTC<fl>
    blockMem[9] = 8'ha;  //JCD<fl><od>
    blockMem[10] = 8'h2b;  //JCA<fl>
    blockMem[11] = 8'hc;  //JCD<fl><od>
    blockMem[12] = 8'h2d;  //JCA<fl>
    blockMem[13] = 8'hf;  //JCD<fl><od>
    blockMem[14] = 8'h33;  //CCD<fl><od>
    blockMem[15] = 8'h3d;  //CCA<fl>
    blockMem[16] = 8'hc;  //JCD<fl><od>
    blockMem[17] = 8'h4e;  //RTC<fl>
    blockMem[18] = 8'h9d;  //SBI<rn><od>
    blockMem[19] = 8'h48;  //RTC<fl>
    blockMem[20] = 8'he;  //JCD<fl><od>
    blockMem[21] = 8'h40;  //INC<rn>
    blockMem[22] = 8'h2a;  //JCA<fl>
    blockMem[23] = 8'h31;  //CCD<fl><od>
    blockMem[24] = 8'h32;  //CCD<fl><od>
    blockMem[25] = 8'h62;  //STA<rn>
    blockMem[26] = 8'h14;  //MVD<rn>
    blockMem[27] = 8'h29;  //JCA<fl>
    blockMem[28] = 8'h48;  //RTC<fl>
    blockMem[29] = 8'h4b;  //RTC<fl>
    blockMem[30] = 8'hf;  //JCD<fl><od>
    blockMem[31] = 8'h30;  //CCD<fl><od>
    blockMem[32] = 8'h8;  //JCD<fl><od>
    blockMem[33] = 8'h33;  //CCD<fl><od>
    blockMem[34] = 8'h3f;  //CCA<fl>
    blockMem[35] = 8'h2a;  //JCA<fl>
    blockMem[36] = 8'hb;  //JCD<fl><od>
    blockMem[37] = 8'h5b;  //MVI<rn><od>
    blockMem[38] = 8'h39;  //CCA<fl>
    blockMem[39] = 8'h2e;  //JCA<fl>
    blockMem[40] = 8'h9;  //JCD<fl><od>
    blockMem[41] = 8'h63;  //STA<rn>
    blockMem[42] = 8'h4d;  //RTC<fl>
    blockMem[43] = 8'h5b;  //MVI<rn><od>
    blockMem[44] = 8'hd;  //JCD<fl><od>
    blockMem[45] = 8'h48;  //RTC<fl>
    blockMem[46] = 8'h66;  //STA<rn>
    blockMem[47] = 8'h11;  //MVD<rn>
    blockMem[48] = 8'h38;  //CCA<fl>
    blockMem[49] = 8'h50;  //DCR<rn>
    blockMem[50] = 8'h80;  //ADA<rn>
    blockMem[51] = 8'h4c;  //RTC<fl>
    blockMem[52] = 8'h7f;  //POP<rn>
    blockMem[53] = 8'ha;  //JCD<fl><od>
    blockMem[54] = 8'h8;  //JCD<fl><od>
    blockMem[55] = 8'h37;  //CCD<fl><od>
    blockMem[56] = 8'h92;  //SBA<rn>
    blockMem[57] = 8'hec;  //XRI<rn><od>
    blockMem[58] = 8'h69;  //PSH<rn>
    blockMem[59] = 8'h45;  //INC<rn>
    blockMem[60] = 8'h2f;  //JCA<fl>
    blockMem[61] = 8'h8;  //JCD<fl><od>
    blockMem[62] = 8'h28;  //JCA<fl>
    blockMem[63] = 8'h78;  //POP<rn>
    blockMem[64] = 8'h73;  //LDA<rn>
    blockMem[65] = 8'h35;  //CCD<fl><od>
    blockMem[66] = 8'h2b;  //JCA<fl>
    blockMem[67] = 8'h18;  //RSP
    blockMem[68] = 8'h2a;  //JCA<fl>
    blockMem[69] = 8'h91;  //SBA<rn>
    blockMem[70] = 8'h48;  //RTC<fl>
    blockMem[71] = 8'h49;  //RTC<fl>
    blockMem[72] = 8'h7c;  //POP<rn>
    blockMem[73] = 8'hdc;  //ORI<rn><od>
    blockMem[74] = 8'h28;  //JCA<fl>
    blockMem[75] = 8'h48;  //RTC<fl>
    blockMem[76] = 8'h3d;  //CCA<fl>
    blockMem[77] = 8'h7b;  //POP<rn>
    blockMem[78] = 8'h6d;  //PSH<rn>
    blockMem[79] = 8'hca;  //ANI<rn><od>
    blockMem[80] = 8'h35;  //CCD<fl><od>
    blockMem[81] = 8'h48;  //RTC<fl>
    blockMem[82] = 8'h31;  //CCD<fl><od>
    blockMem[83] = 8'h4e;  //RTC<fl>
    blockMem[84] = 8'h2d;  //JCA<fl>
    blockMem[85] = 8'h3d;  //CCA<fl>
    blockMem[86] = 8'h3d;  //CCA<fl>
    blockMem[87] = 8'h57;  //DCR<rn>
    blockMem[88] = 8'hc;  //JCD<fl><od>
    blockMem[89] = 8'h4c;  //RTC<fl>
    blockMem[90] = 8'h35;  //CCD<fl><od>
    blockMem[91] = 8'h28;  //JCA<fl>
    blockMem[92] = 8'h6f;  //PSH<rn>
    blockMem[93] = 8'h37;  //CCD<fl><od>
    blockMem[94] = 8'h2c;  //JCA<fl>
    blockMem[95] = 8'h38;  //CCA<fl>
    blockMem[96] = 8'h49;  //RTC<fl>
    blockMem[97] = 8'hc;  //JCD<fl><od>
    blockMem[98] = 8'h36;  //CCD<fl><od>
    blockMem[99] = 8'ha2;  //ACA<rn>
    blockMem[100] = 8'h44;  //INC<rn>
    blockMem[101] = 8'hf;  //JCD<fl><od>
    blockMem[102] = 8'h8d;  //ADI<rn><od>
    blockMem[103] = 8'h4f;  //RTC<fl>
    blockMem[104] = 8'h2e;  //JCA<fl>
    blockMem[105] = 8'h1f;  //MVS<rn>
    blockMem[106] = 8'h2c;  //JCA<fl>
    blockMem[107] = 8'h4f;  //RTC<fl>
    blockMem[108] = 8'hd;  //JCD<fl><od>
    blockMem[109] = 8'hbf;  //SCI<rn><od>
    blockMem[110] = 8'hc;  //JCD<fl><od>
    blockMem[111] = 8'h55;  //DCR<rn>
    blockMem[112] = 8'h2e;  //JCA<fl>
    blockMem[113] = 8'h17;  //MVD<rn>
    blockMem[114] = 8'hf;  //JCD<fl><od>
    blockMem[115] = 8'h5c;  //MVI<rn><od>
    blockMem[116] = 8'h6e;  //PSH<rn>
    blockMem[117] = 8'h33;  //CCD<fl><od>
    blockMem[118] = 8'h29;  //JCA<fl>
    blockMem[119] = 8'hdb;  //ORI<rn><od>
    blockMem[120] = 8'h65;  //STA<rn>
    blockMem[121] = 8'h4c;  //RTC<fl>
    blockMem[122] = 8'h16;  //MVD<rn>
    blockMem[123] = 8'hb;  //JCD<fl><od>
    blockMem[124] = 8'h5a;  //MVI<rn><od>
    blockMem[125] = 8'h35;  //CCD<fl><od>
    blockMem[126] = 8'h63;  //STA<rn>
    blockMem[127] = 8'h72;  //LDA<rn>
    blockMem[128] = 8'h3f;  //CCA<fl>
    blockMem[129] = 8'ha;  //JCD<fl><od>
    blockMem[130] = 8'h16;  //MVD<rn>
    blockMem[131] = 8'h4b;  //RTC<fl>
    blockMem[132] = 8'he;  //JCD<fl><od>
    blockMem[133] = 8'h96;  //SBA<rn>
    blockMem[134] = 8'h4d;  //RTC<fl>
    blockMem[135] = 8'hbd;  //SCI<rn><od>
    blockMem[136] = 8'h3c;  //CCA<fl>
    blockMem[137] = 8'h2f;  //JCA<fl>
    blockMem[138] = 8'hdb;  //ORI<rn><od>
    blockMem[139] = 8'h5a;  //MVI<rn><od>
    blockMem[140] = 8'h34;  //CCD<fl><od>
    blockMem[141] = 8'h77;  //LDA<rn>
    blockMem[142] = 8'hf;  //JCD<fl><od>
    blockMem[143] = 8'hae;  //ACI<rn><od>
    blockMem[144] = 8'h36;  //CCD<fl><od>
    blockMem[145] = 8'h5a;  //MVI<rn><od>
    blockMem[146] = 8'h64;  //STA<rn>
    blockMem[147] = 8'h4b;  //RTC<fl>
    blockMem[148] = 8'h3b;  //CCA<fl>
    blockMem[149] = 8'h5e;  //MVI<rn><od>
    blockMem[150] = 8'h2a;  //JCA<fl>
    blockMem[151] = 8'h2c;  //JCA<fl>
    blockMem[152] = 8'h30;  //CCD<fl><od>
    blockMem[153] = 8'h2e;  //JCA<fl>
    blockMem[154] = 8'h53;  //DCR<rn>
    blockMem[155] = 8'h19;  //MVS<rn>
    blockMem[156] = 8'hc;  //JCD<fl><od>
    blockMem[157] = 8'h8a;  //ADI<rn><od>
    blockMem[158] = 8'hd4;  //ORA<rn>
    blockMem[159] = 8'h3d;  //CCA<fl>
    blockMem[160] = 8'hc9;  //ANI<rn><od>
    blockMem[161] = 8'ha7;  //ACA<rn>
    blockMem[162] = 8'h33;  //CCD<fl><od>
    blockMem[163] = 8'hf;  //JCD<fl><od>
    blockMem[164] = 8'h3b;  //CCA<fl>
    blockMem[165] = 8'h77;  //LDA<rn>
    blockMem[166] = 8'h49;  //RTC<fl>
    blockMem[167] = 8'h39;  //CCA<fl>
    blockMem[168] = 8'h10;  //LSP
    blockMem[169] = 8'h37;  //CCD<fl><od>
    blockMem[170] = 8'h33;  //CCD<fl><od>
    blockMem[171] = 8'hb9;  //SCI<rn><od>
    blockMem[172] = 8'h9;  //JCD<fl><od>
    blockMem[173] = 8'h10;  //LSP
    blockMem[174] = 8'h5f;  //MVI<rn><od>
    blockMem[175] = 8'hc;  //JCD<fl><od>
    blockMem[176] = 8'h50;  //DCR<rn>
    blockMem[177] = 8'h3c;  //CCA<fl>
    blockMem[178] = 8'h35;  //CCD<fl><od>
    blockMem[179] = 8'hb9;  //SCI<rn><od>
    blockMem[180] = 8'h34;  //CCD<fl><od>
    blockMem[181] = 8'he5;  //XRA<rn>
    blockMem[182] = 8'h2c;  //JCA<fl>
    blockMem[183] = 8'h4b;  //RTC<fl>
    blockMem[184] = 8'h49;  //RTC<fl>
    blockMem[185] = 8'h4b;  //RTC<fl>
    blockMem[186] = 8'had;  //ACI<rn><od>
    blockMem[187] = 8'h3e;  //CCA<fl>
    blockMem[188] = 8'h61;  //STA<rn>
    blockMem[189] = 8'h3d;  //CCA<fl>
    blockMem[190] = 8'h49;  //RTC<fl>
    blockMem[191] = 8'hb;  //JCD<fl><od>
    blockMem[192] = 8'h69;  //PSH<rn>
    blockMem[193] = 8'hcd;  //ANI<rn><od>
    blockMem[194] = 8'h30;  //CCD<fl><od>
    blockMem[195] = 8'he9;  //XRI<rn><od>
    blockMem[196] = 8'h8b;  //ADI<rn><od>
    blockMem[197] = 8'h39;  //CCA<fl>
    blockMem[198] = 8'h4b;  //RTC<fl>
    blockMem[199] = 8'h68;  //PSH<rn>
    blockMem[200] = 8'h68;  //PSH<rn>
    blockMem[201] = 8'h4d;  //RTC<fl>
    blockMem[202] = 8'h52;  //DCR<rn>
    blockMem[203] = 8'h2d;  //JCA<fl>
    blockMem[204] = 8'hae;  //ACI<rn><od>
    blockMem[205] = 8'hee;  //XRI<rn><od>
    blockMem[206] = 8'h7d;  //POP<rn>
    blockMem[207] = 8'h6a;  //PSH<rn>
    blockMem[208] = 8'h9e;  //SBI<rn><od>
    blockMem[209] = 8'h4e;  //RTC<fl>
    blockMem[210] = 8'h38;  //CCA<fl>
    blockMem[211] = 8'h30;  //CCD<fl><od>
    blockMem[212] = 8'h6b;  //PSH<rn>
    blockMem[213] = 8'h37;  //CCD<fl><od>
    blockMem[214] = 8'he5;  //XRA<rn>
    blockMem[215] = 8'h2e;  //JCA<fl>
    blockMem[216] = 8'ha6;  //ACA<rn>
    blockMem[217] = 8'ha;  //JCD<fl><od>
    blockMem[218] = 8'h4f;  //RTC<fl>
    blockMem[219] = 8'h81;  //ADA<rn>
    blockMem[220] = 8'h39;  //CCA<fl>
    blockMem[221] = 8'hbb;  //SCI<rn><od>
    blockMem[222] = 8'h2a;  //JCA<fl>
    blockMem[223] = 8'h31;  //CCD<fl><od>
    blockMem[224] = 8'h82;  //ADA<rn>
    blockMem[225] = 8'h2d;  //JCA<fl>
    blockMem[226] = 8'h32;  //CCD<fl><od>
    blockMem[227] = 8'haa;  //ACI<rn><od>
    blockMem[228] = 8'h76;  //LDA<rn>
    blockMem[229] = 8'h2c;  //JCA<fl>
    blockMem[230] = 8'h1f;  //MVS<rn>
    blockMem[231] = 8'h5a;  //MVI<rn><od>
    blockMem[232] = 8'hea;  //XRI<rn><od>
    blockMem[233] = 8'h3e;  //CCA<fl>
    blockMem[234] = 8'hc8;  //ANI<rn><od>
    blockMem[235] = 8'h67;  //STA<rn>
    blockMem[236] = 8'h4b;  //RTC<fl>
    blockMem[237] = 8'h30;  //CCD<fl><od>
    blockMem[238] = 8'h30;  //CCD<fl><od>
    blockMem[239] = 8'ha;  //JCD<fl><od>
    blockMem[240] = 8'h69;  //PSH<rn>
    blockMem[241] = 8'h33;  //CCD<fl><od>
    blockMem[242] = 8'h3f;  //CCA<fl>
    blockMem[243] = 8'hec;  //XRI<rn><od>
    blockMem[244] = 8'h38;  //CCA<fl>
    blockMem[245] = 8'h4f;  //RTC<fl>
    blockMem[246] = 8'ha4;  //ACA<rn>
    blockMem[247] = 8'h78;  //POP<rn>
    blockMem[248] = 8'h4d;  //RTC<fl>
    blockMem[249] = 8'h5c;  //MVI<rn><od>
    blockMem[250] = 8'h79;  //POP<rn>
    blockMem[251] = 8'hce;  //ANI<rn><od>
    blockMem[252] = 8'h3d;  //CCA<fl>
    blockMem[253] = 8'hba;  //SCI<rn><od>
    blockMem[254] = 8'h3b;  //CCA<fl>
    blockMem[255] = 8'h4c;  //RTC<fl
    *//*
    blockMem[0] = 8'h01; //CLR
    blockMem[1] = 8'h2e;  //JCA<fl>
    blockMem[2] = 8'ha6;  //ACA<rn>
    blockMem[3] = 8'h8;  //JCD<fl><od>
    blockMem[4] = 8'h49;  //RTC<fl>
    blockMem[5] = 8'h39;  //CCA<fl>
    blockMem[6] = 8'h2e;  //JCA<fl>
    blockMem[7] = 8'h3a;  //CCA<fl>
    blockMem[8] = 8'h7b;  //POP<rn>
    blockMem[9] = 8'hd6;  //ORA<rn>
    blockMem[10] = 8'h4c;  //RTC<fl>
    blockMem[11] = 8'he6;  //XRA<rn>
    blockMem[12] = 8'h75;  //LDA<rn>
    blockMem[13] = 8'hf;  //JCD<fl><od>
    blockMem[14] = 8'h2c;  //JCA<fl>
    blockMem[15] = 8'h5f;  //MVI<rn><od>
    blockMem[16] = 8'h49;  //RTC<fl>
    blockMem[17] = 8'h4b;  //RTC<fl>
    blockMem[18] = 8'h2e;  //JCA<fl>
    blockMem[19] = 8'hc;  //JCD<fl><od>
    blockMem[20] = 8'h17;  //MVD<rn>
    blockMem[21] = 8'h65;  //STA<rn>
    blockMem[22] = 8'h4c;  //RTC<fl>
    blockMem[23] = 8'h34;  //CCD<fl><od>
    blockMem[24] = 8'h80;  //ADA<rn>
    blockMem[25] = 8'hbc;  //SCI<rn><od>
    blockMem[26] = 8'he;  //JCD<fl><od>
    blockMem[27] = 8'ha;  //JCD<fl><od>
    blockMem[28] = 8'hf;  //JCD<fl><od>
    blockMem[29] = 8'h49;  //RTC<fl>
    blockMem[30] = 8'hb2;  //SCA<rn>
    blockMem[31] = 8'h3d;  //CCA<fl>
    blockMem[32] = 8'h19;  //MVS<rn>
    blockMem[33] = 8'h4d;  //RTC<fl>
    blockMem[34] = 8'h3e;  //CCA<fl>
    blockMem[35] = 8'h4b;  //RTC<fl>
    blockMem[36] = 8'h48;  //RTC<fl>
    blockMem[37] = 8'h3e;  //CCA<fl>
    blockMem[38] = 8'he;  //JCD<fl><od>
    blockMem[39] = 8'h4b;  //RTC<fl>
    blockMem[40] = 8'h10;  //LSP
    blockMem[41] = 8'h29;  //JCA<fl>
    blockMem[42] = 8'hc6;  //ANA<rn>
    blockMem[43] = 8'h1f;  //MVS<rn>
    blockMem[44] = 8'h97;  //SBA<rn>
    blockMem[45] = 8'h26;  //NOT<rn>
    blockMem[46] = 8'hd4;  //ORA<rn>
    blockMem[47] = 8'h46;  //INC<rn>
    blockMem[48] = 8'hbc;  //SCI<rn><od>
    blockMem[49] = 8'hb;  //JCD<fl><od>
    blockMem[50] = 8'h4a;  //RTC<fl>
    blockMem[51] = 8'hab;  //ACI<rn><od>
    blockMem[52] = 8'h9;  //JCD<fl><od>
    blockMem[53] = 8'h8;  //JCD<fl><od>
    blockMem[54] = 8'h4e;  //RTC<fl>
    blockMem[55] = 8'h78;  //POP<rn>
    blockMem[56] = 8'h28;  //JCA<fl>
    blockMem[57] = 8'h37;  //CCD<fl><od>
    blockMem[58] = 8'h21;  //NOT<rn>
    blockMem[59] = 8'hb0;  //SCA<rn>
    blockMem[60] = 8'h48;  //RTC<fl>
    blockMem[61] = 8'h2b;  //JCA<fl>
    blockMem[62] = 8'hc;  //JCD<fl><od>
    blockMem[63] = 8'hd5;  //ORA<rn>
    blockMem[64] = 8'h6f;  //PSH<rn>
    blockMem[65] = 8'h2d;  //JCA<fl>
    blockMem[66] = 8'h4a;  //RTC<fl>
    blockMem[67] = 8'h12;  //MVD<rn>
    blockMem[68] = 8'h9d;  //SBI<rn><od>
    blockMem[69] = 8'h3e;  //CCA<fl>
    blockMem[70] = 8'he5;  //XRA<rn>
    blockMem[71] = 8'h71;  //LDA<rn>
    blockMem[72] = 8'h38;  //CCA<fl>
    blockMem[73] = 8'h39;  //CCA<fl>
    blockMem[74] = 8'hf;  //JCD<fl><od>
    blockMem[75] = 8'h10;  //LSP
    blockMem[76] = 8'h18;  //RSP
    blockMem[77] = 8'h24;  //NOT<rn>
    blockMem[78] = 8'hd9;  //ORI<rn><od>
    blockMem[79] = 8'ha0;  //ACA<rn>
    blockMem[80] = 8'h5e;  //MVI<rn><od>
    blockMem[81] = 8'h3e;  //CCA<fl>
    blockMem[82] = 8'h1c;  //MVS<rn>
    blockMem[83] = 8'h2b;  //JCA<fl>
    blockMem[84] = 8'ha;  //JCD<fl><od>
    blockMem[85] = 8'h73;  //LDA<rn>
    blockMem[86] = 8'h13;  //MVD<rn>
    blockMem[87] = 8'h4a;  //RTC<fl>
    blockMem[88] = 8'h80;  //ADA<rn>
    blockMem[89] = 8'h89;  //ADI<rn><od>
    blockMem[90] = 8'h49;  //RTC<fl>
    blockMem[91] = 8'ha7;  //ACA<rn>
    blockMem[92] = 8'h4d;  //RTC<fl>
    blockMem[93] = 8'h3b;  //CCA<fl>
    blockMem[94] = 8'h5b;  //MVI<rn><od>
    blockMem[95] = 8'h65;  //STA<rn>
    blockMem[96] = 8'h26;  //NOT<rn>
    blockMem[97] = 8'hea;  //XRI<rn><od>
    blockMem[98] = 8'ha;  //JCD<fl><od>
    blockMem[99] = 8'h2d;  //JCA<fl>
    blockMem[100] = 8'ha;  //JCD<fl><od>
    blockMem[101] = 8'hc;  //JCD<fl><od>
    blockMem[102] = 8'h48;  //RTC<fl>
    blockMem[103] = 8'h67;  //STA<rn>
    blockMem[104] = 8'h2f;  //JCA<fl>
    blockMem[105] = 8'hdd;  //ORI<rn><od>
    blockMem[106] = 8'h67;  //STA<rn>
    blockMem[107] = 8'h5b;  //MVI<rn><od>
    blockMem[108] = 8'hc;  //JCD<fl><od>
    blockMem[109] = 8'h4d;  //RTC<fl>
    blockMem[110] = 8'h4a;  //RTC<fl>
    blockMem[111] = 8'h1a;  //MVS<rn>
    blockMem[112] = 8'h5a;  //MVI<rn><od>
    blockMem[113] = 8'hb3;  //SCA<rn>
    blockMem[114] = 8'h4a;  //RTC<fl>
    blockMem[115] = 8'h3a;  //CCA<fl>
    blockMem[116] = 8'h10;  //LSP
    blockMem[117] = 8'h69;  //PSH<rn>
    blockMem[118] = 8'h8b;  //ADI<rn><od>
    blockMem[119] = 8'h2;  //CLC
    blockMem[120] = 8'h64;  //STA<rn>
    blockMem[121] = 8'h3e;  //CCA<fl>
    blockMem[122] = 8'h8c;  //ADI<rn><od>
    blockMem[123] = 8'h7b;  //POP<rn>
    blockMem[124] = 8'h37;  //CCD<fl><od>
    blockMem[125] = 8'h34;  //CCD<fl><od>
    blockMem[126] = 8'h49;  //RTC<fl>
    blockMem[127] = 8'h83;  //ADA<rn>
    blockMem[128] = 8'h38;  //CCA<fl>
    blockMem[129] = 8'had;  //ACI<rn><od>
    blockMem[130] = 8'h49;  //RTC<fl>
    blockMem[131] = 8'h71;  //LDA<rn>
    blockMem[132] = 8'h76;  //LDA<rn>
    blockMem[133] = 8'h3d;  //CCA<fl>
    blockMem[134] = 8'h4e;  //RTC<fl>
    blockMem[135] = 8'h12;  //MVD<rn>
    blockMem[136] = 8'h3b;  //CCA<fl>
    blockMem[137] = 8'h3b;  //CCA<fl>
    blockMem[138] = 8'h61;  //STA<rn>
    blockMem[139] = 8'h35;  //CCD<fl><od>
    blockMem[140] = 8'h11;  //MVD<rn>
    blockMem[141] = 8'h43;  //INC<rn>
    blockMem[142] = 8'h86;  //ADA<rn>
    blockMem[143] = 8'hb6;  //SCA<rn>
    blockMem[144] = 8'hf;  //JCD<fl><od>
    blockMem[145] = 8'h5b;  //MVI<rn><od>
    blockMem[146] = 8'hc8;  //ANI<rn><od>
    blockMem[147] = 8'h8;  //JCD<fl><od>
    blockMem[148] = 8'h1c;  //MVS<rn>
    blockMem[149] = 8'h2e;  //JCA<fl>
    blockMem[150] = 8'h3f;  //CCA<fl>
    blockMem[151] = 8'h5f;  //MVI<rn><od>
    blockMem[152] = 8'h3f;  //CCA<fl>
    blockMem[153] = 8'h37;  //CCD<fl><od>
    blockMem[154] = 8'h3c;  //CCA<fl>
    blockMem[155] = 8'h94;  //SBA<rn>
    blockMem[156] = 8'h1a;  //MVS<rn>
    blockMem[157] = 8'h2f;  //JCA<fl>
    blockMem[158] = 8'h2f;  //JCA<fl>
    blockMem[159] = 8'h27;  //NOT<rn>
    blockMem[160] = 8'h67;  //STA<rn>
    blockMem[161] = 8'hba;  //SCI<rn><od>
    blockMem[162] = 8'hf;  //JCD<fl><od>
    blockMem[163] = 8'ha5;  //ACA<rn>
    blockMem[164] = 8'h36;  //CCD<fl><od>
    blockMem[165] = 8'h3a;  //CCA<fl>
    blockMem[166] = 8'h33;  //CCD<fl><od>
    blockMem[167] = 8'hc;  //JCD<fl><od>
    blockMem[168] = 8'h78;  //POP<rn>
    blockMem[169] = 8'hdf;  //ORI<rn><od>
    blockMem[170] = 8'h39;  //CCA<fl>
    blockMem[171] = 8'h9;  //JCD<fl><od>
    blockMem[172] = 8'h1f;  //MVS<rn>
    blockMem[173] = 8'hb1;  //SCA<rn>
    blockMem[174] = 8'hba;  //SCI<rn><od>
    blockMem[175] = 8'h7b;  //POP<rn>
    blockMem[176] = 8'h29;  //JCA<fl>
    blockMem[177] = 8'hd;  //JCD<fl><od>
    blockMem[178] = 8'h9;  //JCD<fl><od>
    blockMem[179] = 8'h8e;  //ADI<rn><od>
    blockMem[180] = 8'h41;  //INC<rn>
    blockMem[181] = 8'h15;  //MVD<rn>
    blockMem[182] = 8'hdc;  //ORI<rn><od>
    blockMem[183] = 8'h3f;  //CCA<fl>
    blockMem[184] = 8'h10;  //LSP
    blockMem[185] = 8'h13;  //MVD<rn>
    blockMem[186] = 8'h5c;  //MVI<rn><od>
    blockMem[187] = 8'hd;  //JCD<fl><od>
    blockMem[188] = 8'he2;  //XRA<rn>
    blockMem[189] = 8'h47;  //INC<rn>
    blockMem[190] = 8'h9b;  //SBI<rn><od>
    blockMem[191] = 8'hd2;  //ORA<rn>
    blockMem[192] = 8'ha;  //JCD<fl><od>
    blockMem[193] = 8'h62;  //STA<rn>
    blockMem[194] = 8'hea;  //XRI<rn><od>
    blockMem[195] = 8'h37;  //CCD<fl><od>
    blockMem[196] = 8'h2e;  //JCA<fl>
    blockMem[197] = 8'h2a;  //JCA<fl>
    blockMem[198] = 8'h2e;  //JCA<fl>
    blockMem[199] = 8'h8a;  //ADI<rn><od>
    blockMem[200] = 8'h7c;  //POP<rn>
    blockMem[201] = 8'h4d;  //RTC<fl>
    blockMem[202] = 8'h2a;  //JCA<fl>
    blockMem[203] = 8'h3e;  //CCA<fl>
    blockMem[204] = 8'h64;  //STA<rn>
    blockMem[205] = 8'h5c;  //MVI<rn><od>
    blockMem[206] = 8'h16;  //MVD<rn>
    blockMem[207] = 8'h36;  //CCD<fl><od>
    blockMem[208] = 8'h12;  //MVD<rn>
    blockMem[209] = 8'hb7;  //SCA<rn>
    blockMem[210] = 8'h35;  //CCD<fl><od>
    blockMem[211] = 8'h20;  //NOT<rn>
    blockMem[212] = 8'h6d;  //PSH<rn>
    blockMem[213] = 8'h33;  //CCD<fl><od>
    blockMem[214] = 8'h6a;  //PSH<rn>
    blockMem[215] = 8'h2b;  //JCA<fl>
    blockMem[216] = 8'hc;  //JCD<fl><od>
    blockMem[217] = 8'h6b;  //PSH<rn>
    blockMem[218] = 8'h91;  //SBA<rn>
    blockMem[219] = 8'h4a;  //RTC<fl>
    blockMem[220] = 8'h29;  //JCA<fl>
    blockMem[221] = 8'ha;  //JCD<fl><od>
    blockMem[222] = 8'h48;  //RTC<fl>
    blockMem[223] = 8'h30;  //CCD<fl><od>
    blockMem[224] = 8'h1e;  //MVS<rn>
    blockMem[225] = 8'h74;  //LDA<rn>
    blockMem[226] = 8'h82;  //ADA<rn>
    blockMem[227] = 8'h78;  //POP<rn>
    blockMem[228] = 8'he8;  //XRI<rn><od>
    blockMem[229] = 8'h33;  //CCD<fl><od>
    blockMem[230] = 8'hf;  //JCD<fl><od>
    blockMem[231] = 8'ha;  //JCD<fl><od>
    blockMem[232] = 8'h13;  //MVD<rn>
    blockMem[233] = 8'h3a;  //CCA<fl>
    blockMem[234] = 8'h2;  //CLC
    blockMem[235] = 8'h23;  //NOT<rn>
    blockMem[236] = 8'h3b;  //CCA<fl>
    blockMem[237] = 8'hed;  //XRI<rn><od>
    blockMem[238] = 8'hd0;  //ORA<rn>
    blockMem[239] = 8'h74;  //LDA<rn>
    blockMem[240] = 8'ha;  //JCD<fl><od>
    blockMem[241] = 8'h9;  //JCD<fl><od>
    blockMem[242] = 8'h19;  //MVS<rn>
    blockMem[243] = 8'h39;  //CCA<fl>
    blockMem[244] = 8'h28;  //JCA<fl>
    blockMem[245] = 8'h49;  //RTC<fl>
    blockMem[246] = 8'ha;  //JCD<fl><od>
    blockMem[247] = 8'h63;  //STA<rn>
    blockMem[248] = 8'h9;  //JCD<fl><od>
    blockMem[249] = 8'h42;  //INC<rn>
    blockMem[250] = 8'ha;  //JCD<fl><od>
    blockMem[251] = 8'h3c;  //CCA<fl>
    blockMem[252] = 8'h37;  //CCD<fl><od>
    blockMem[253] = 8'h6e;  //PSH<rn>
    blockMem[254] = 8'h84;  //ADA<rn>
    blockMem[255] = 8'h65;  //STA<rn>
    */
    /*blockMem[0] = 8'h01;  //SBA<rn>
    blockMem[1] = 8'h40;  //JCA<fl>
    blockMem[2] = 8'hc9;  //ANI<rn><od>
    blockMem[3] = 8'h6d;  //PSH<rn>
    blockMem[4] = 8'ha3;  //ACA<rn>
    blockMem[5] = 8'h7b;  //POP<rn>
    blockMem[6] = 8'hd8;  //ORI<rn><od>
    blockMem[7] = 8'h75;  //LDA<rn>
    blockMem[8] = 8'ha7;  //ACA<rn>
    blockMem[9] = 8'h1a;  //MVS<rn>
    blockMem[10] = 8'h6f;  //PSH<rn>
    blockMem[11] = 8'h3d;  //CCA<fl>
    blockMem[12] = 8'h51;  //DCR<rn>
    blockMem[13] = 8'h5d;  //MVI<rn><od>
    blockMem[14] = 8'h69;  //PSH<rn>
    blockMem[15] = 8'h1a;  //MVS<rn>
    blockMem[16] = 8'h7f;  //POP<rn>
    blockMem[17] = 8'hd8;  //ORI<rn><od>
    blockMem[18] = 8'h6d;  //PSH<rn>
    blockMem[19] = 8'h45;  //INC<rn>
    blockMem[20] = 8'h30;  //CCD<fl><od>
    blockMem[21] = 8'h1b;  //MVS<rn>
    blockMem[22] = 8'h8d;  //ADI<rn><od>
    blockMem[23] = 8'h2c;  //JCA<fl>
    blockMem[24] = 8'h68;  //PSH<rn>
    blockMem[25] = 8'h78;  //POP<rn>
    blockMem[26] = 8'h19;  //MVS<rn>
    blockMem[27] = 8'h5e;  //MVI<rn><od>
    blockMem[28] = 8'hb7;  //SCA<rn>
    blockMem[29] = 8'hc3;  //ANA<rn>
    blockMem[30] = 8'h18;  //RSP
    blockMem[31] = 8'haa;  //ACI<rn><od>
    blockMem[32] = 8'h13;  //MVD<rn>
    blockMem[33] = 8'h76;  //LDA<rn>
    blockMem[34] = 8'h3d;  //CCA<fl>
    blockMem[35] = 8'h1d;  //MVS<rn>
    blockMem[36] = 8'hc0;  //ANA<rn>
    blockMem[37] = 8'h63;  //STA<rn>
    blockMem[38] = 8'h5c;  //MVI<rn><od>
    blockMem[39] = 8'heb;  //XRI<rn><od>
    blockMem[40] = 8'hd9;  //ORI<rn><od>
    blockMem[41] = 8'hc8;  //ANI<rn><od>
    blockMem[42] = 8'h1f;  //MVS<rn>
    blockMem[43] = 8'h8b;  //ADI<rn><od>
    blockMem[44] = 8'h34;  //CCD<fl><od>
    blockMem[45] = 8'h92;  //SBA<rn>
    blockMem[46] = 8'he1;  //XRA<rn>
    blockMem[47] = 8'haa;  //ACI<rn><od>
    blockMem[48] = 8'hd;  //JCD<fl><od>
    blockMem[49] = 8'hc9;  //ANI<rn><od>
    blockMem[50] = 8'h7a;  //POP<rn>
    blockMem[51] = 8'h1e;  //MVS<rn>
    blockMem[52] = 8'he6;  //XRA<rn>
    blockMem[53] = 8'ha5;  //ACA<rn>
    blockMem[54] = 8'h1c;  //MVS<rn>
    blockMem[55] = 8'h67;  //STA<rn>
    blockMem[56] = 8'h35;  //CCD<fl><od>
    blockMem[57] = 8'h6f;  //PSH<rn>
    blockMem[58] = 8'h43;  //INC<rn>
    blockMem[59] = 8'h77;  //LDA<rn>
    blockMem[60] = 8'h1e;  //MVS<rn>
    blockMem[61] = 8'h5d;  //MVI<rn><od>
    blockMem[62] = 8'hcb;  //ANI<rn><od>
    blockMem[63] = 8'h63;  //STA<rn>
    blockMem[64] = 8'h7f;  //POP<rn>
    blockMem[65] = 8'h18;  //RSP
    blockMem[66] = 8'h76;  //LDA<rn>
    blockMem[67] = 8'he5;  //XRA<rn>
    blockMem[68] = 8'h84;  //ADA<rn>
    blockMem[69] = 8'h7e;  //POP<rn>
    blockMem[70] = 8'h2d;  //JCA<fl>
    blockMem[71] = 8'h5b;  //MVI<rn><od>
    blockMem[72] = 8'hcf;  //ANI<rn><od>
    blockMem[73] = 8'h65;  //STA<rn>
    blockMem[74] = 8'h6f;  //PSH<rn>
    blockMem[75] = 8'hcc;  //ANI<rn><od>
    blockMem[76] = 8'h56;  //DCR<rn>
    blockMem[77] = 8'h23;  //NOT<rn>
    blockMem[78] = 8'ha7;  //ACA<rn>
    blockMem[79] = 8'hcf;  //ANI<rn><od>
    blockMem[80] = 8'h84;  //ADA<rn>
    blockMem[81] = 8'h13;  //MVD<rn>
    blockMem[82] = 8'h6b;  //PSH<rn>
    blockMem[83] = 8'h3a;  //CCA<fl>
    blockMem[84] = 8'h5d;  //MVI<rn><od>
    blockMem[85] = 8'h85;  //ADA<rn>
    blockMem[86] = 8'ha;  //JCD<fl><od>
    blockMem[87] = 8'h5b;  //MVI<rn><od>
    blockMem[88] = 8'h98;  //SBI<rn><od>
    blockMem[89] = 8'h1d;  //MVS<rn>
    blockMem[90] = 8'h58;  //MVI<rn><od>
    blockMem[91] = 8'h79;  //POP<rn>
    blockMem[92] = 8'h19;  //MVS<rn>
    blockMem[93] = 8'h79;  //POP<rn>
    blockMem[94] = 8'h69;  //PSH<rn>
    blockMem[95] = 8'h33;  //CCD<fl><od>
    blockMem[96] = 8'h91;  //SBA<rn>
    blockMem[97] = 8'h5c;  //MVI<rn><od>
    blockMem[98] = 8'hdf;  //ORI<rn><od>
    blockMem[99] = 8'h1a;  //MVS<rn>
    blockMem[100] = 8'h36;  //CCD<fl><od>
    blockMem[101] = 8'h22;  //NOT<rn>
    blockMem[102] = 8'h7a;  //POP<rn>
    blockMem[103] = 8'h55;  //DCR<rn>
    blockMem[104] = 8'h60;  //RLA
    blockMem[105] = 8'h6d;  //PSH<rn>
    blockMem[106] = 8'h3c;  //CCA<fl>
    blockMem[107] = 8'h1b;  //MVS<rn>
    blockMem[108] = 8'hc;  //JCD<fl><od>
    blockMem[109] = 8'h36;  //CCD<fl><od>
    blockMem[110] = 8'h14;  //MVD<rn>
    blockMem[111] = 8'h6f;  //PSH<rn>
    blockMem[112] = 8'h97;  //SBA<rn>
    blockMem[113] = 8'hb0;  //SCA<rn>
    blockMem[114] = 8'h6e;  //PSH<rn>
    blockMem[115] = 8'h5d;  //MVI<rn><od>
    blockMem[116] = 8'h6d;  //PSH<rn>
    blockMem[117] = 8'h5e;  //MVI<rn><od>
    blockMem[118] = 8'h2e;  //JCA<fl>
    blockMem[119] = 8'h69;  //PSH<rn>
    blockMem[120] = 8'h75;  //LDA<rn>
    blockMem[121] = 8'h67;  //STA<rn>
    blockMem[122] = 8'he1;  //XRA<rn>
    blockMem[123] = 8'h97;  //SBA<rn>
    blockMem[124] = 8'h11;  //MVD<rn>
    blockMem[125] = 8'h91;  //SBA<rn>
    blockMem[126] = 8'h5f;  //MVI<rn><od>
    blockMem[127] = 8'h3f;  //CCA<fl>
    blockMem[128] = 8'he4;  //XRA<rn>
    blockMem[129] = 8'h48;  //RTC<fl>
    blockMem[130] = 8'h42;  //INC<rn>
    blockMem[131] = 8'h46;  //INC<rn>
    blockMem[132] = 8'h85;  //ADA<rn>
    blockMem[133] = 8'h7f;  //POP<rn>
    blockMem[134] = 8'h61;  //STA<rn>
    blockMem[135] = 8'h56;  //DCR<rn>
    blockMem[136] = 8'h7c;  //POP<rn>
    blockMem[137] = 8'hb7;  //SCA<rn>
    blockMem[138] = 8'h72;  //LDA<rn>
    blockMem[139] = 8'h71;  //LDA<rn>
    blockMem[140] = 8'h9f;  //SBI<rn><od>
    blockMem[141] = 8'h1c;  //MVS<rn>
    blockMem[142] = 8'he7;  //XRA<rn>
    blockMem[143] = 8'h46;  //INC<rn>
    blockMem[144] = 8'h76;  //LDA<rn>
    blockMem[145] = 8'h12;  //MVD<rn>
    blockMem[146] = 8'h50;  //DCR<rn>
    blockMem[147] = 8'h73;  //LDA<rn>
    blockMem[148] = 8'h7b;  //POP<rn>
    blockMem[149] = 8'h9d;  //SBI<rn><od>
    blockMem[150] = 8'h7d;  //POP<rn>
    blockMem[151] = 8'hb1;  //SCA<rn>
    blockMem[152] = 8'h22;  //NOT<rn>
    blockMem[153] = 8'hb5;  //SCA<rn>
    blockMem[154] = 8'h51;  //DCR<rn>
    blockMem[155] = 8'h45;  //INC<rn>
    blockMem[156] = 8'hcc;  //ANI<rn><od>
    blockMem[157] = 8'h9a;  //SBI<rn><od>
    blockMem[158] = 8'hbb;  //SCI<rn><od>
    blockMem[159] = 8'h29;  //JCA<fl>
    blockMem[160] = 8'h37;  //CCD<fl><od>
    blockMem[161] = 8'h3e;  //CCA<fl>
    blockMem[162] = 8'h5c;  //MVI<rn><od>
    blockMem[163] = 8'hed;  //XRI<rn><od>
    blockMem[164] = 8'h15;  //MVD<rn>
    blockMem[165] = 8'h18;  //RSP
    blockMem[166] = 8'h1d;  //MVS<rn>
    blockMem[167] = 8'h9d;  //SBI<rn><od>
    blockMem[168] = 8'h73;  //LDA<rn>
    blockMem[169] = 8'he1;  //XRA<rn>
    blockMem[170] = 8'h72;  //LDA<rn>
    blockMem[171] = 8'hc7;  //ANA<rn>
    blockMem[172] = 8'h13;  //MVD<rn>
    blockMem[173] = 8'h90;  //SBA<rn>
    blockMem[174] = 8'h19;  //MVS<rn>
    blockMem[175] = 8'h4a;  //RTC<fl>
    blockMem[176] = 8'h38;  //CCA<fl>
    blockMem[177] = 8'h9d;  //SBI<rn><od>
    blockMem[178] = 8'h1d;  //MVS<rn>
    blockMem[179] = 8'h7d;  //POP<rn>
    blockMem[180] = 8'h22;  //NOT<rn>
    blockMem[181] = 8'h1d;  //MVS<rn>
    blockMem[182] = 8'ha5;  //ACA<rn>
    blockMem[183] = 8'h7e;  //POP<rn>
    blockMem[184] = 8'h86;  //ADA<rn>
    blockMem[185] = 8'h1c;  //MVS<rn>
    blockMem[186] = 8'hd1;  //ORA<rn>
    blockMem[187] = 8'h7e;  //POP<rn>
    blockMem[188] = 8'hc7;  //ANA<rn>
    blockMem[189] = 8'hb7;  //SCA<rn>
    blockMem[190] = 8'h9d;  //SBI<rn><od>
    blockMem[191] = 8'h79;  //POP<rn>
    blockMem[192] = 8'hea;  //XRI<rn><od>
    blockMem[193] = 8'h1e;  //MVS<rn>
    blockMem[194] = 8'ha5;  //ACA<rn>
    blockMem[195] = 8'h1d;  //MVS<rn>
    blockMem[196] = 8'h64;  //STA<rn>
    blockMem[197] = 8'h13;  //MVD<rn>
    blockMem[198] = 8'h7e;  //POP<rn>
    blockMem[199] = 8'ha3;  //ACA<rn>
    blockMem[200] = 8'h12;  //MVD<rn>
    blockMem[201] = 8'h55;  //DCR<rn>
    blockMem[202] = 8'h59;  //MVI<rn><od>
    blockMem[203] = 8'h72;  //LDA<rn>
    blockMem[204] = 8'h7d;  //POP<rn>
    blockMem[205] = 8'h17;  //MVD<rn>
    blockMem[206] = 8'h47;  //INC<rn>
    blockMem[207] = 8'hd1;  //ORA<rn>
    blockMem[208] = 8'h2c;  //JCA<fl>
    blockMem[209] = 8'he1;  //XRA<rn>
    blockMem[210] = 8'h6d;  //PSH<rn>
    blockMem[211] = 8'h2b;  //JCA<fl>
    blockMem[212] = 8'h2a;  //JCA<fl>
    blockMem[213] = 8'h6b;  //PSH<rn>
    blockMem[214] = 8'hcc;  //ANI<rn><od>
    blockMem[215] = 8'h3e;  //CCA<fl>
    blockMem[216] = 8'h7e;  //POP<rn>
    blockMem[217] = 8'h79;  //POP<rn>
    blockMem[218] = 8'h2a;  //JCA<fl>
    blockMem[219] = 8'hbb;  //SCI<rn><od>
    blockMem[220] = 8'h7a;  //POP<rn>
    blockMem[221] = 8'hc3;  //ANA<rn>
    blockMem[222] = 8'hab;  //ACI<rn><od>
    blockMem[223] = 8'h6d;  //PSH<rn>
    blockMem[224] = 8'h55;  //DCR<rn>
    blockMem[225] = 8'h65;  //STA<rn>
    blockMem[226] = 8'h6f;  //PSH<rn>
    blockMem[227] = 8'ha;  //JCD<fl><od>
    blockMem[228] = 8'hcd;  //ANI<rn><od>
    blockMem[229] = 8'hb2;  //SCA<rn>
    blockMem[230] = 8'h2;  //CLC
    blockMem[231] = 8'haf;  //ACI<rn><od>
    blockMem[232] = 8'h69;  //PSH<rn>
    blockMem[233] = 8'h97;  //SBA<rn>
    blockMem[234] = 8'h75;  //LDA<rn>
    blockMem[235] = 8'hb1;  //SCA<rn>
    blockMem[236] = 8'hc;  //JCD<fl><od>
    blockMem[237] = 8'h18;  //RSP
    blockMem[238] = 8'h48;  //RTC<fl>
    blockMem[239] = 8'hde;  //ORI<rn><od>
    blockMem[240] = 8'h64;  //STA<rn>
    blockMem[241] = 8'h98;  //SBI<rn><od>
    blockMem[242] = 8'h85;  //ADA<rn>
    blockMem[243] = 8'h63;  //STA<rn>
    blockMem[244] = 8'h6b;  //PSH<rn>
    blockMem[245] = 8'h2f;  //JCA<fl>
    blockMem[246] = 8'h4b;  //RTC<fl>
    blockMem[247] = 8'hc;  //JCD<fl><od>
    blockMem[248] = 8'hc0;  //ANA<rn>
    blockMem[249] = 8'h3f;  //CCA<fl>
    blockMem[250] = 8'h9c;  //SBI<rn><od>
    blockMem[251] = 8'hcf;  //ANI<rn><od>
    blockMem[252] = 8'h1;  //CLR
    blockMem[253] = 8'h15;  //MVD<rn>
    blockMem[254] = 8'h7c;  //POP<rn>
    blockMem[255] = 8'h01; //CLR
<<<<<<< HEAD
    */  /*  
        blockMem[0] = 8'h01;  //CLR
=======
    */    
        /*blockMem[0] = 8'h01;  //CLR
>>>>>>> e083d40d6961653dcdb4f46b0cb8c2cea20102bd
        blockMem[1] = 8'h1f;  //MVS<rn>
        blockMem[2] = 8'h62;  //STA<rn>
        blockMem[3] = 8'h9c;  //SBI<rn><od>
        blockMem[4] = 8'h54;  //DCR<rn>
        blockMem[5] = 8'he5;  //XRA<rn>
        blockMem[6] = 8'hb2;  //SCA<rn>
        blockMem[7] = 8'h62;  //STA<rn>
        blockMem[8] = 8'hb6;  //SCA<rn>
        blockMem[9] = 8'h47;  //INC<rn>
        blockMem[10] = 8'h58;  //MVI<rn><od>
        blockMem[11] = 8'h5b;  //MVI<rn><od>
        blockMem[12] = 8'he4;  //XRA<rn>
        blockMem[13] = 8'hb6;  //SCA<rn>
        blockMem[14] = 8'h7d;  //POP<rn>
        blockMem[15] = 8'h7b;  //POP<rn>
        blockMem[16] = 8'h61;  //STA<rn>
        blockMem[17] = 8'h79;  //POP<rn>
        blockMem[18] = 8'h5e;  //MVI<rn><od>
        blockMem[19] = 8'h13;  //MVD<rn>
        blockMem[20] = 8'h86;  //ADA<rn>
        blockMem[21] = 8'h83;  //ADA<rn>
        blockMem[22] = 8'h58;  //MVI<rn><od>
        blockMem[23] = 8'hed;  //XRI<rn><od>
        blockMem[24] = 8'h6f;  //PSH<rn>
        blockMem[25] = 8'hcc;  //ANI<rn><od>
        blockMem[26] = 8'h18;  //RSP
        blockMem[27] = 8'hea;  //XRI<rn><od>
        blockMem[28] = 8'h5a;  //MVI<rn><od>
        blockMem[29] = 8'h59;  //MVI<rn><od>
        blockMem[30] = 8'h1f;  //MVS<rn>
        blockMem[31] = 8'h00;  //SBA<rn>
        blockMem[32] = 8'hdd;  //ORI<rn><od>
        blockMem[33] = 8'h22;  //NOT<rn>
        blockMem[34] = 8'h6c;  //PSH<rn>
        blockMem[35] = 8'h6d;  //PSH<rn>
        blockMem[36] = 8'h62;  //STA<rn>
        blockMem[37] = 8'h5e;  //MVI<rn><od>
        blockMem[38] = 8'h8d;  //ADI<rn><od>
        blockMem[39] = 8'h9b;  //SBI<rn><od>
        blockMem[40] = 8'h11;  //MVD<rn>
        blockMem[41] = 8'h00;  //ACA<rn>
        blockMem[42] = 8'h76;  //LDA<rn>
        blockMem[43] = 8'he6;  //XRA<rn>
        blockMem[44] = 8'h77;  //LDA<rn>
        blockMem[45] = 8'h71;  //LDA<rn>
        blockMem[46] = 8'hd9;  //ORI<rn><od>
        blockMem[47] = 8'h17;  //MVD<rn>
        blockMem[48] = 8'h67;  //STA<rn>
        blockMem[49] = 8'h97;  //SBA<rn>
        blockMem[50] = 8'h24;  //NOT<rn>
        blockMem[51] = 8'h19;  //MVS<rn>
        blockMem[52] = 8'h71;  //LDA<rn>
        blockMem[53] = 8'h61;  //STA<rn>
        blockMem[54] = 8'h6c;  //PSH<rn>
        blockMem[55] = 8'h61;  //STA<rn>
        blockMem[56] = 8'h1a;  //MVS<rn>
        blockMem[57] = 8'ha3;  //ACA<rn>
        blockMem[58] = 8'hdb;  //ORI<rn><od>
        blockMem[59] = 8'h13;  //MVD<rn>
        blockMem[60] = 8'h58;  //MVI<rn><od>
        blockMem[61] = 8'h68;  //PSH<rn>
        blockMem[62] = 8'h14;  //MVD<rn>
        blockMem[63] = 8'hbe;  //SCI<rn><od>
        blockMem[64] = 8'hc8;  //ANI<rn><od>
        blockMem[65] = 8'h6a;  //PSH<rn>
        blockMem[66] = 8'h57;  //DCR<rn>
        blockMem[67] = 8'h22;  //NOT<rn>
        blockMem[68] = 8'h67;  //STA<rn>
        blockMem[69] = 8'haf;  //ACI<rn><od>
        blockMem[70] = 8'h5c;  //MVI<rn><od>
        blockMem[71] = 8'h5d;  //MVI<rn><od>
        blockMem[72] = 8'h6f;  //PSH<rn>
        blockMem[73] = 8'h6c;  //PSH<rn>
        blockMem[74] = 8'hbb;  //SCI<rn><od>
        blockMem[75] = 8'h7d;  //POP<rn>
        blockMem[76] = 8'hd8;  //ORI<rn><od>
        blockMem[77] = 8'h68;  //PSH<rn>
        blockMem[78] = 8'h7c;  //POP<rn>
        blockMem[79] = 8'h77;  //LDA<rn>
        blockMem[80] = 8'h58;  //MVI<rn><od>
        blockMem[81] = 8'h7f;  //POP<rn>
        blockMem[82] = 8'h13;  //MVD<rn>
        blockMem[83] = 8'hde;  //ORI<rn><od>
        blockMem[84] = 8'h71;  //LDA<rn>
        blockMem[85] = 8'h8e;  //ADI<rn><od>
        blockMem[86] = 8'h42;  //INC<rn>
        blockMem[87] = 8'h6a;  //PSH<rn>
        blockMem[88] = 8'ha5;  //ACA<rn>
        blockMem[89] = 8'hd6;  //ORA<rn>
        blockMem[90] = 8'h11;  //MVD<rn>
        blockMem[91] = 8'h63;  //STA<rn>
        blockMem[92] = 8'hd2;  //ORA<rn>
        blockMem[93] = 8'hc3;  //ANA<rn>
        blockMem[94] = 8'h11;  //MVD<rn>
        blockMem[95] = 8'h62;  //STA<rn>
        blockMem[96] = 8'hb4;  //SCA<rn>
        blockMem[97] = 8'h66;  //STA<rn>
        blockMem[98] = 8'hd0;  //ORA<rn>
        blockMem[99] = 8'h6a;  //PSH<rn>
        blockMem[100] = 8'h69;  //PSH<rn>
        blockMem[101] = 8'h1d;  //MVS<rn>
        blockMem[102] = 8'ha2;  //ACA<rn>
        blockMem[103] = 8'heb;  //XRI<rn><od>
        blockMem[104] = 8'h54;  //DCR<rn>
        blockMem[105] = 8'h19;  //MVS<rn>
        blockMem[106] = 8'h5a;  //MVI<rn><od>
        blockMem[107] = 8'hbc;  //SCI<rn><od>
        blockMem[108] = 8'h93;  //SBA<rn>
        blockMem[109] = 8'he8;  //XRI<rn><od>
        blockMem[110] = 8'h69;  //PSH<rn>
        blockMem[111] = 8'h99;  //SBI<rn><od>
        blockMem[112] = 8'h7d;  //POP<rn>
        blockMem[113] = 8'ha7;  //ACA<rn>
        blockMem[114] = 8'h26;  //NOT<rn>
        blockMem[115] = 8'h91;  //SBA<rn>
        blockMem[116] = 8'hbe;  //SCI<rn><od>
        blockMem[117] = 8'h6a;  //PSH<rn>
        blockMem[118] = 8'hd5;  //ORA<rn>
        blockMem[119] = 8'hc4;  //ANA<rn>
        blockMem[120] = 8'h66;  //STA<rn>
        blockMem[121] = 8'h79;  //POP<rn>
        blockMem[122] = 8'h61;  //STA<rn>
        blockMem[123] = 8'hb2;  //SCA<rn>
        blockMem[124] = 8'hc3;  //ANA<rn>
        blockMem[125] = 8'h7e;  //POP<rn>
        blockMem[126] = 8'h6d;  //PSH<rn>
        blockMem[127] = 8'h97;  //SBA<rn>
        blockMem[128] = 8'h6f;  //PSH<rn>
        blockMem[129] = 8'haa;  //ACI<rn><od>
        blockMem[130] = 8'h00;  //ACA<rn>
        blockMem[131] = 8'h61;  //STA<rn>
        blockMem[132] = 8'h96;  //SBA<rn>
        blockMem[133] = 8'he9;  //XRI<rn><od>
        blockMem[134] = 8'h65;  //STA<rn>
        blockMem[135] = 8'h61;  //STA<rn>
        blockMem[136] = 8'h10;  //LSP
        blockMem[137] = 8'h7d;  //POP<rn>
        blockMem[138] = 8'h17;  //MVD<rn>
        blockMem[139] = 8'h58;  //MVI<rn><od>
        blockMem[140] = 8'h66;  //STA<rn>
        blockMem[141] = 8'h7a;  //POP<rn>
        blockMem[142] = 8'h79;  //POP<rn>
        blockMem[143] = 8'h7b;  //POP<rn>
        blockMem[144] = 8'h11;  //MVD<rn>
        blockMem[145] = 8'h69;  //PSH<rn>
        blockMem[146] = 8'hd3;  //ORA<rn>
        blockMem[147] = 8'h7f;  //POP<rn>
        blockMem[148] = 8'h20;  //NOT<rn>
        blockMem[149] = 8'h6a;  //PSH<rn>
        blockMem[150] = 8'h7a;  //POP<rn>
        blockMem[151] = 8'h5c;  //MVI<rn><od>
        blockMem[152] = 8'h27;  //NOT<rn>
        blockMem[153] = 8'h1c;  //MVS<rn>
        blockMem[154] = 8'h6f;  //PSH<rn>
        blockMem[155] = 8'h61;  //STA<rn>
        blockMem[156] = 8'hc3;  //ANA<rn>
        blockMem[157] = 8'hef;  //XRI<rn><od>
        blockMem[158] = 8'h68;  //PSH<rn>
        blockMem[159] = 8'h78;  //POP<rn>
        blockMem[160] = 8'h40;  //INC<rn>
        blockMem[161] = 8'h98;  //SBI<rn><od>
        blockMem[162] = 8'h6a;  //PSH<rn>
        blockMem[163] = 8'h7d;  //POP<rn>
        blockMem[164] = 8'h65;  //STA<rn>
        blockMem[165] = 8'h1d;  //MVS<rn>
        blockMem[166] = 8'hbf;  //SCI<rn><od>
        blockMem[167] = 8'h6b;  //PSH<rn>
        blockMem[168] = 8'h73;  //LDA<rn>
        blockMem[169] = 8'h55;  //DCR<rn>
        blockMem[170] = 8'hbb;  //SCI<rn><od>
        blockMem[171] = 8'hc2;  //ANA<rn>
        blockMem[172] = 8'h73;  //LDA<rn>
        blockMem[173] = 8'hd3;  //ORA<rn>
        blockMem[174] = 8'h58;  //MVI<rn><od>
        blockMem[175] = 8'h67;  //STA<rn>
        blockMem[176] = 8'h5d;  //MVI<rn><od>
        blockMem[177] = 8'h25;  //NOT<rn>
        blockMem[178] = 8'h5e;  //MVI<rn><od>
        blockMem[179] = 8'h40;  //INC<rn>
        blockMem[180] = 8'h7c;  //POP<rn>
        blockMem[181] = 8'h1f;  //MVS<rn>
        blockMem[182] = 8'h6e;  //PSH<rn>
        blockMem[183] = 8'hdf;  //ORI<rn><od>
        blockMem[184] = 8'hce;  //ANI<rn><od>
        blockMem[185] = 8'h63;  //STA<rn>
        blockMem[186] = 8'h5d;  //MVI<rn><od>
        blockMem[187] = 8'hcc;  //ANI<rn><od>
        blockMem[188] = 8'h5d;  //MVI<rn><od>
        blockMem[189] = 8'h43;  //INC<rn>
        blockMem[190] = 8'h51;  //DCR<rn>
        blockMem[191] = 8'h76;  //LDA<rn>
        blockMem[192] = 8'h6f;  //PSH<rn>
        blockMem[193] = 8'h14;  //MVD<rn>
        blockMem[194] = 8'h59;  //MVI<rn><od>
        blockMem[195] = 8'h62;  //STA<rn>
        blockMem[196] = 8'hde;  //ORI<rn><od>
        blockMem[197] = 8'h51;  //DCR<rn>
        blockMem[198] = 8'h5e;  //MVI<rn><od>
        blockMem[199] = 8'h6a;  //PSH<rn>
        blockMem[200] = 8'h62;  //STA<rn>
        blockMem[201] = 8'h73;  //LDA<rn>
        blockMem[202] = 8'h69;  //PSH<rn>
        blockMem[203] = 8'h7a;  //POP<rn>
        blockMem[204] = 8'h64;  //STA<rn>
        blockMem[205] = 8'h76;  //LDA<rn>
        blockMem[206] = 8'h1b;  //MVS<rn>
        blockMem[207] = 8'h58;  //MVI<rn><od>
        blockMem[208] = 8'h69;  //PSH<rn>
        blockMem[209] = 8'h78;  //POP<rn>
        blockMem[210] = 8'h1a;  //MVS<rn>
        blockMem[211] = 8'h9e;  //SBI<rn><od>
        blockMem[212] = 8'h94;  //SBA<rn>
        blockMem[213] = 8'h78;  //POP<rn>
        blockMem[214] = 8'h92;  //SBA<rn>
        blockMem[215] = 8'h65;  //STA<rn>
        blockMem[216] = 8'h20;  //NOT<rn>
        blockMem[217] = 8'h7a;  //POP<rn>
        blockMem[218] = 8'h77;  //LDA<rn>
        blockMem[219] = 8'h2;  //CLC
        blockMem[220] = 8'h59;  //MVI<rn><od>
        blockMem[221] = 8'h77;  //LDA<rn>
        blockMem[222] = 8'h5b;  //MVI<rn><od>
        blockMem[223] = 8'h00;  //ACA<rn>
        blockMem[224] = 8'h66;  //STA<rn>
        blockMem[225] = 8'h8a;  //ADI<rn><od>
        blockMem[226] = 8'h17;  //MVD<rn>
        blockMem[227] = 8'hec;  //XRI<rn><od>
        blockMem[228] = 8'h5d;  //MVI<rn><od>
        blockMem[229] = 8'h59;  //MVI<rn><od>
        blockMem[230] = 8'he7;  //XRA<rn>
        blockMem[231] = 8'h1a;  //MVS<rn>
        blockMem[232] = 8'h74;  //LDA<rn>
        blockMem[233] = 8'h5d;  //MVI<rn><od>
        blockMem[234] = 8'h88;  //ADI<rn><od>
        blockMem[235] = 8'h1b;  //MVS<rn>
        blockMem[236] = 8'h15;  //MVD<rn>
        blockMem[237] = 8'h67;  //STA<rn>
        blockMem[238] = 8'h77;  //LDA<rn>
        blockMem[239] = 8'h42;  //INC<rn>
        blockMem[240] = 8'he1;  //XRA<rn>
        blockMem[241] = 8'h66;  //STA<rn>
        blockMem[242] = 8'hbe;  //SCI<rn><od>
        blockMem[243] = 8'h41;  //INC<rn>
        blockMem[244] = 8'hce;  //ANI<rn><od>
        blockMem[245] = 8'h45;  //INC<rn>
        blockMem[246] = 8'h7f;  //POP<rn>
        blockMem[247] = 8'h88;  //ADI<rn><od>
        blockMem[248] = 8'h53;  //DCR<rn>
        blockMem[249] = 8'h79;  //POP<rn>
        blockMem[250] = 8'h6d;  //PSH<rn>
        blockMem[251] = 8'h62;  //STA<rn>
        blockMem[252] = 8'h9a;  //SBI<rn><od>
        blockMem[253] = 8'hef;  //XRI<rn><od>
        blockMem[254] = 8'h7c;  //POP<rn>
        blockMem[255] = 8'h01;  //CLR
*/
blockMem[0] = 8'h01;  //SBA<rn>
blockMem[1] = 8'h58;  //JCA<fl>
blockMem[2] = 8'hc9;  //ANI<rn><od>
blockMem[3] = 8'h6d;  //PSH<rn>
blockMem[4] = 8'ha3;  //ACA<rn>
blockMem[5] = 8'h7b;  //POP<rn>
blockMem[6] = 8'hd8;  //ORI<rn><od>
blockMem[7] = 8'h75;  //LDA<rn>
blockMem[8] = 8'ha7;  //ACA<rn>
blockMem[9] = 8'h1a;  //MVS<rn>
blockMem[10] = 8'h6f;  //PSH<rn>
blockMem[11] = 8'h3d;  //CCA<fl>
blockMem[12] = 8'h51;  //DCR<rn>
blockMem[13] = 8'h5d;  //MVI<rn><od>
blockMem[14] = 8'h69;  //PSH<rn>
blockMem[15] = 8'h1a;  //MVS<rn>
blockMem[16] = 8'h7f;  //POP<rn>
blockMem[17] = 8'hd8;  //ORI<rn><od>
blockMem[18] = 8'h6d;  //PSH<rn>
blockMem[19] = 8'h45;  //INC<rn>
blockMem[20] = 8'h30;  //CCD<fl><od>
blockMem[21] = 8'h1b;  //MVS<rn>
blockMem[22] = 8'h8d;  //ADI<rn><od>
blockMem[23] = 8'h2c;  //JCA<fl>
blockMem[24] = 8'h68;  //PSH<rn>
blockMem[25] = 8'h78;  //POP<rn>
blockMem[26] = 8'h19;  //MVS<rn>
blockMem[27] = 8'h5e;  //MVI<rn><od>
blockMem[28] = 8'hb7;  //SCA<rn>
blockMem[29] = 8'hc3;  //ANA<rn>
blockMem[30] = 8'h18;  //RSP
blockMem[31] = 8'haa;  //ACI<rn><od>
blockMem[32] = 8'h13;  //MVD<rn>
blockMem[33] = 8'h76;  //LDA<rn>
blockMem[34] = 8'h3d;  //CCA<fl>
blockMem[35] = 8'h1d;  //MVS<rn>
blockMem[36] = 8'hc0;  //ANA<rn>
blockMem[37] = 8'h63;  //STA<rn>
blockMem[38] = 8'h5c;  //MVI<rn><od>
blockMem[39] = 8'heb;  //XRI<rn><od>
blockMem[40] = 8'hd9;  //ORI<rn><od>
blockMem[41] = 8'hc8;  //ANI<rn><od>
blockMem[42] = 8'h1f;  //MVS<rn>
blockMem[43] = 8'h8b;  //ADI<rn><od>
blockMem[44] = 8'h34;  //CCD<fl><od>
blockMem[45] = 8'h92;  //SBA<rn>
blockMem[46] = 8'he1;  //XRA<rn>
blockMem[47] = 8'haa;  //ACI<rn><od>
blockMem[48] = 8'hd;  //JCD<fl><od>
blockMem[49] = 8'hc9;  //ANI<rn><od>
blockMem[50] = 8'h7a;  //POP<rn>
blockMem[51] = 8'h1e;  //MVS<rn>
blockMem[52] = 8'he6;  //XRA<rn>
blockMem[53] = 8'ha5;  //ACA<rn>
blockMem[54] = 8'h1c;  //MVS<rn>
blockMem[55] = 8'h67;  //STA<rn>
blockMem[56] = 8'h35;  //CCD<fl><od>
blockMem[57] = 8'h6f;  //PSH<rn>
blockMem[58] = 8'h43;  //INC<rn>
blockMem[59] = 8'h77;  //LDA<rn>
blockMem[60] = 8'h1e;  //MVS<rn>
blockMem[61] = 8'h5d;  //MVI<rn><od>
blockMem[62] = 8'hcb;  //ANI<rn><od>
blockMem[63] = 8'h63;  //STA<rn>
blockMem[64] = 8'h7f;  //POP<rn>
blockMem[65] = 8'h18;  //RSP
blockMem[66] = 8'h76;  //LDA<rn>
blockMem[67] = 8'he5;  //XRA<rn>
blockMem[68] = 8'h84;  //ADA<rn>
blockMem[69] = 8'h7e;  //POP<rn>
blockMem[70] = 8'h2d;  //JCA<fl>
blockMem[71] = 8'h5b;  //MVI<rn><od>
blockMem[72] = 8'hcf;  //ANI<rn><od>
blockMem[73] = 8'h65;  //STA<rn>
blockMem[74] = 8'h6f;  //PSH<rn>
blockMem[75] = 8'hcc;  //ANI<rn><od>
blockMem[76] = 8'h56;  //DCR<rn>
blockMem[77] = 8'h23;  //NOT<rn>
blockMem[78] = 8'ha7;  //ACA<rn>
blockMem[79] = 8'hcf;  //ANI<rn><od>
blockMem[80] = 8'h84;  //ADA<rn>
blockMem[81] = 8'h13;  //MVD<rn>
blockMem[82] = 8'h6b;  //PSH<rn>
blockMem[83] = 8'h3a;  //CCA<fl>
blockMem[84] = 8'h5d;  //MVI<rn><od>
blockMem[85] = 8'h85;  //ADA<rn>
blockMem[86] = 8'ha;  //JCD<fl><od>
blockMem[87] = 8'h5b;  //MVI<rn><od>
blockMem[88] = 8'h98;  //SBI<rn><od>
blockMem[89] = 8'h1d;  //MVS<rn>
blockMem[90] = 8'h58;  //MVI<rn><od>
blockMem[91] = 8'h79;  //POP<rn>
blockMem[92] = 8'h19;  //MVS<rn>
blockMem[93] = 8'h79;  //POP<rn>
blockMem[94] = 8'h69;  //PSH<rn>
blockMem[95] = 8'h33;  //CCD<fl><od>
blockMem[96] = 8'h91;  //SBA<rn>
blockMem[97] = 8'h5c;  //MVI<rn><od>
blockMem[98] = 8'hdf;  //ORI<rn><od>
blockMem[99] = 8'h1a;  //MVS<rn>
blockMem[100] = 8'h36;  //CCD<fl><od>
blockMem[101] = 8'h22;  //NOT<rn>
blockMem[102] = 8'h7a;  //POP<rn>
blockMem[103] = 8'h55;  //DCR<rn>
blockMem[104] = 8'h60;  //RLA
blockMem[105] = 8'h6d;  //PSH<rn>
blockMem[106] = 8'h3c;  //CCA<fl>
blockMem[107] = 8'h1b;  //MVS<rn>
blockMem[108] = 8'hc;  //JCD<fl><od>
blockMem[109] = 8'h36;  //CCD<fl><od>
blockMem[110] = 8'h14;  //MVD<rn>
blockMem[111] = 8'h6f;  //PSH<rn>
blockMem[112] = 8'h97;  //SBA<rn>
blockMem[113] = 8'hb0;  //SCA<rn>
blockMem[114] = 8'h6e;  //PSH<rn>
blockMem[115] = 8'h5d;  //MVI<rn><od>
blockMem[116] = 8'h6d;  //PSH<rn>
blockMem[117] = 8'h5e;  //MVI<rn><od>
blockMem[118] = 8'h2e;  //JCA<fl>
blockMem[119] = 8'h69;  //PSH<rn>
blockMem[120] = 8'h75;  //LDA<rn>
blockMem[121] = 8'h67;  //STA<rn>
blockMem[122] = 8'he1;  //XRA<rn>
blockMem[123] = 8'h97;  //SBA<rn>
blockMem[124] = 8'h11;  //MVD<rn>
blockMem[125] = 8'h91;  //SBA<rn>
blockMem[126] = 8'h5f;  //MVI<rn><od>
blockMem[127] = 8'h3f;  //CCA<fl>
blockMem[128] = 8'he4;  //XRA<rn>
blockMem[129] = 8'h48;  //RTC<fl>
blockMem[130] = 8'h42;  //INC<rn>
blockMem[131] = 8'h46;  //INC<rn>
blockMem[132] = 8'h85;  //ADA<rn>
blockMem[133] = 8'h7f;  //POP<rn>
blockMem[134] = 8'h61;  //STA<rn>
blockMem[135] = 8'h56;  //DCR<rn>
blockMem[136] = 8'h7c;  //POP<rn>
blockMem[137] = 8'hb7;  //SCA<rn>
blockMem[138] = 8'h72;  //LDA<rn>
blockMem[139] = 8'h71;  //LDA<rn>
blockMem[140] = 8'h9f;  //SBI<rn><od>
blockMem[141] = 8'h1c;  //MVS<rn>
blockMem[142] = 8'he7;  //XRA<rn>
blockMem[143] = 8'h46;  //INC<rn>
blockMem[144] = 8'h76;  //LDA<rn>
blockMem[145] = 8'h12;  //MVD<rn>
blockMem[146] = 8'h50;  //DCR<rn>
blockMem[147] = 8'h73;  //LDA<rn>
blockMem[148] = 8'h7b;  //POP<rn>
blockMem[149] = 8'h9d;  //SBI<rn><od>
blockMem[150] = 8'h7d;  //POP<rn>
blockMem[151] = 8'hb1;  //SCA<rn>
blockMem[152] = 8'h22;  //NOT<rn>
blockMem[153] = 8'hb5;  //SCA<rn>
blockMem[154] = 8'h51;  //DCR<rn>
blockMem[155] = 8'h45;  //INC<rn>
blockMem[156] = 8'hcc;  //ANI<rn><od>
blockMem[157] = 8'h9a;  //SBI<rn><od>
blockMem[158] = 8'hbb;  //SCI<rn><od>
blockMem[159] = 8'h29;  //JCA<fl>
blockMem[160] = 8'h37;  //CCD<fl><od>
blockMem[161] = 8'h3e;  //CCA<fl>
blockMem[162] = 8'h5c;  //MVI<rn><od>
blockMem[163] = 8'hed;  //XRI<rn><od>
blockMem[164] = 8'h15;  //MVD<rn>
blockMem[165] = 8'h18;  //RSP
blockMem[166] = 8'h1d;  //MVS<rn>
blockMem[167] = 8'h9d;  //SBI<rn><od>
blockMem[168] = 8'h73;  //LDA<rn>
blockMem[169] = 8'he1;  //XRA<rn>
blockMem[170] = 8'h72;  //LDA<rn>
blockMem[171] = 8'hc7;  //ANA<rn>
blockMem[172] = 8'h13;  //MVD<rn>
blockMem[173] = 8'h90;  //SBA<rn>
blockMem[174] = 8'h19;  //MVS<rn>
blockMem[175] = 8'h4a;  //RTC<fl>
blockMem[176] = 8'h38;  //CCA<fl>
blockMem[177] = 8'h9d;  //SBI<rn><od>
blockMem[178] = 8'h1d;  //MVS<rn>
blockMem[179] = 8'h7d;  //POP<rn>
blockMem[180] = 8'h22;  //NOT<rn>
blockMem[181] = 8'h1d;  //MVS<rn>
blockMem[182] = 8'ha5;  //ACA<rn>
blockMem[183] = 8'h7e;  //POP<rn>
blockMem[184] = 8'h86;  //ADA<rn>
blockMem[185] = 8'h1c;  //MVS<rn>
blockMem[186] = 8'hd1;  //ORA<rn>
blockMem[187] = 8'h7e;  //POP<rn>
blockMem[188] = 8'hc7;  //ANA<rn>
blockMem[189] = 8'hb7;  //SCA<rn>
blockMem[190] = 8'h9d;  //SBI<rn><od>
blockMem[191] = 8'h79;  //POP<rn>
blockMem[192] = 8'hea;  //XRI<rn><od>
blockMem[193] = 8'h1e;  //MVS<rn>
blockMem[194] = 8'ha5;  //ACA<rn>
blockMem[195] = 8'h1d;  //MVS<rn>
blockMem[196] = 8'h64;  //STA<rn>
blockMem[197] = 8'h13;  //MVD<rn>
blockMem[198] = 8'h7e;  //POP<rn>
blockMem[199] = 8'ha3;  //ACA<rn>
blockMem[200] = 8'h12;  //MVD<rn>
blockMem[201] = 8'h55;  //DCR<rn>
blockMem[202] = 8'h59;  //MVI<rn><od>
blockMem[203] = 8'h72;  //LDA<rn>
blockMem[204] = 8'h7d;  //POP<rn>
blockMem[205] = 8'h17;  //MVD<rn>
blockMem[206] = 8'h47;  //INC<rn>
blockMem[207] = 8'hd1;  //ORA<rn>
blockMem[208] = 8'h2c;  //JCA<fl>
blockMem[209] = 8'he1;  //XRA<rn>
blockMem[210] = 8'h6d;  //PSH<rn>
blockMem[211] = 8'h2b;  //JCA<fl>
blockMem[212] = 8'h2a;  //JCA<fl>
blockMem[213] = 8'h6b;  //PSH<rn>
blockMem[214] = 8'hcc;  //ANI<rn><od>
blockMem[215] = 8'h3e;  //CCA<fl>
blockMem[216] = 8'h7e;  //POP<rn>
blockMem[217] = 8'h79;  //POP<rn>
blockMem[218] = 8'h2a;  //JCA<fl>
blockMem[219] = 8'hbb;  //SCI<rn><od>
blockMem[220] = 8'h7a;  //POP<rn>
blockMem[221] = 8'hc3;  //ANA<rn>
blockMem[222] = 8'hab;  //ACI<rn><od>
blockMem[223] = 8'h6d;  //PSH<rn>
blockMem[224] = 8'h55;  //DCR<rn>
blockMem[225] = 8'h65;  //STA<rn>
blockMem[226] = 8'h6f;  //PSH<rn>
blockMem[227] = 8'ha;  //JCD<fl><od>
blockMem[228] = 8'hcd;  //ANI<rn><od>
blockMem[229] = 8'hb2;  //SCA<rn>
blockMem[230] = 8'h2;  //CLC
blockMem[231] = 8'haf;  //ACI<rn><od>
blockMem[232] = 8'h69;  //PSH<rn>
blockMem[233] = 8'h97;  //SBA<rn>
blockMem[234] = 8'h75;  //LDA<rn>
blockMem[235] = 8'hb1;  //SCA<rn>
blockMem[236] = 8'hc;  //JCD<fl><od>
blockMem[237] = 8'h18;  //RSP
blockMem[238] = 8'h48;  //RTC<fl>
blockMem[239] = 8'hde;  //ORI<rn><od>
blockMem[240] = 8'h64;  //STA<rn>
blockMem[241] = 8'h98;  //SBI<rn><od>
blockMem[242] = 8'h85;  //ADA<rn>
blockMem[243] = 8'h63;  //STA<rn>
blockMem[244] = 8'h6b;  //PSH<rn>
blockMem[245] = 8'h2f;  //JCA<fl>
blockMem[246] = 8'h4b;  //RTC<fl>
blockMem[247] = 8'hc;  //JCD<fl><od>
blockMem[248] = 8'hc0;  //ANA<rn>
blockMem[249] = 8'h3f;  //CCA<fl>
blockMem[250] = 8'h9c;  //SBI<rn><od>
blockMem[251] = 8'hcf;  //ANI<rn><od>
blockMem[252] = 8'h1;  //CLR
blockMem[253] = 8'h15;  //MVD<rn>
blockMem[254] = 8'h7c;  //POP<rn>
blockMem[255] = 8'h01; //CLR
    /*
         blockMem[0]  = 8'h01;
         blockMem[1]  = 8'h43;
         blockMem[2]  = 8'h0b;
         blockMem[3]  = 8'h01;
         blockMem[4]  = 8'h02;
         blockMem[5]  = 8'h42;
         blockMem[6]  = 8'h0b;
         blockMem[7]  = 8'h01;
         blockMem[8]  = 8'h02;
         blockMem[9]  = 8'h41;
         blockMem[10] = 8'h0b;
         blockMem[11] = 8'h01;
         blockMem[12] = 8'h02;
         blockMem[13] = 8'h40;
         blockMem[14] = 8'hf8;
         blockMem[15] = 8'h0b;
         blockMem[16] = 8'h01;
         blockMem[17] = 8'h00;
         blockMem[18] = 8'h00;
         blockMem[19] = 8'h00;
         blockMem[20] = 8'h00;
         blockMem[21] = 8'h00;
         blockMem[22] = 8'h00;
         blockMem[23] = 8'h00;
         blockMem[24] = 8'h00;
         blockMem[25] = 8'h00;
         blockMem[26] = 8'h00;
         blockMem[27] = 8'h00;
         blockMem[28] = 8'h00;
         blockMem[29] = 8'h00;
         blockMem[30] = 8'h00;
         blockMem[31] = 8'h00;
         blockMem[32] = 8'h00;
         blockMem[33] = 8'h00;
         blockMem[34] = 8'h00;
         blockMem[35] = 8'h00;
         blockMem[36] = 8'h00;
         blockMem[37] = 8'h00;
         blockMem[38] = 8'h00;
         blockMem[39] = 8'h00;
         blockMem[40] = 8'h28;
         blockMem[41] = 8'h29;
         blockMem[42] = 8'h2a;
         blockMem[43] = 8'h2b;
         blockMem[44] = 8'h2c;
         blockMem[45] = 8'h2d;
         blockMem[46] = 8'h2e;
         blockMem[47] = 8'h2f;
         blockMem[48] = 8'h00;
         blockMem[49] = 8'h00;
         blockMem[50] = 8'h00;
         blockMem[51] = 8'h00;
         blockMem[52] = 8'h00;
         blockMem[53] = 8'h00;
         blockMem[54] = 8'h00;
         blockMem[55] = 8'h00;
         blockMem[56] = 8'h00;
         blockMem[57] = 8'h00;
         blockMem[58] = 8'h00;
         blockMem[59] = 8'h00;
         blockMem[60] = 8'h00;
         blockMem[61] = 8'h00;
         blockMem[62] = 8'h00;
         blockMem[63] = 8'h00;
         blockMem[64] = 8'h00;
         blockMem[65] = 8'h00;
         blockMem[66] = 8'h00;
         blockMem[67] = 8'h00;
         blockMem[68] = 8'h00;
         blockMem[69] = 8'h00;
         blockMem[70] = 8'h00;
         blockMem[71] = 8'h00;
         blockMem[72] = 8'h00;
         blockMem[73] = 8'h00;
         blockMem[74] = 8'h00;
         blockMem[75] = 8'h00;
         blockMem[76] = 8'h00;
         blockMem[77] = 8'h00;
         blockMem[78] = 8'h00;
         blockMem[79] = 8'h00;
         blockMem[80] = 8'h00;
         blockMem[81] = 8'h00;
         blockMem[82] = 8'h00;
         blockMem[83] = 8'h00;
         blockMem[84] = 8'h00;
         blockMem[85] = 8'h00;
         blockMem[86] = 8'h00;
         blockMem[87] = 8'h00;
         blockMem[88] = 8'h00;
         blockMem[89] = 8'h00;
         blockMem[90] = 8'h00;
         blockMem[91] = 8'h00;
         blockMem[92] = 8'h00;
         blockMem[93] = 8'h00;
         blockMem[94] = 8'h00;
         blockMem[95] = 8'h00;
         blockMem[96] = 8'h00;
         blockMem[97] = 8'h00;
         blockMem[98] = 8'h00;
         blockMem[99] = 8'h00;
         blockMem[100] =8'h00;
         blockMem[101] =8'h00;
         blockMem[102] =8'h00;
         blockMem[103] =8'h00;
         blockMem[104] =8'h00;
         blockMem[105] =8'h00;
         blockMem[106] =8'h00;
         blockMem[107] =8'h00;
         blockMem[108] =8'h00;
         blockMem[109] =8'h00;
         blockMem[110] =8'h00;
         blockMem[111] =8'h00;
         blockMem[112] =8'h00;
         blockMem[113] =8'h00;
         blockMem[114] =8'h00;
         blockMem[115] =8'h00;
         blockMem[116] =8'h00;
         blockMem[117] =8'h00;
         blockMem[118] =8'h00;
         blockMem[119] =8'h00;
         blockMem[120] =8'h00;
         blockMem[121] =8'h00;
         blockMem[122] =8'h00;
         blockMem[123] =8'h00;
         blockMem[124] =8'h00;
         blockMem[125] =8'h00;
         blockMem[126] =8'h00;
         blockMem[127] =8'h00;
         blockMem[128] =8'h00;
         blockMem[129] =8'h00;
         blockMem[130] =8'h00;
         blockMem[131] =8'h00;
         blockMem[132] =8'h00;
         blockMem[133] =8'h00;
         blockMem[134] =8'h00;
         blockMem[135] =8'h00;
         blockMem[136] =8'h00;
         blockMem[137] =8'h00;
         blockMem[138] =8'h00;
         blockMem[139] =8'h00;
         blockMem[140] =8'h00;
         blockMem[141] =8'h00;
         blockMem[142] =8'h00;
         blockMem[143] =8'h00;
         blockMem[144] =8'h00;
         blockMem[145] =8'h00;
         blockMem[146] =8'h00;
         blockMem[147] =8'h00;
         blockMem[148] =8'h00;
         blockMem[149] =8'h00;
         blockMem[150] =8'h00;
         blockMem[151] =8'h00;
         blockMem[152] =8'h00;
         blockMem[153] =8'h00;
         blockMem[154] =8'h00;
         blockMem[155] =8'h00;
         blockMem[156] =8'h00;
         blockMem[157] =8'h00;
         blockMem[158] =8'h00;
         blockMem[159] =8'h00;
         blockMem[160] =8'h00;
         blockMem[161] =8'h00;
         blockMem[162] =8'h00;
         blockMem[163] =8'h00;
         blockMem[164] =8'h00;
         blockMem[165] =8'h00;
         blockMem[166] =8'h00;
         blockMem[167] =8'h00;
         blockMem[168] =8'h00;
         blockMem[169] =8'h00;
         blockMem[170] =8'h00;
         blockMem[171] =8'h00;
         blockMem[172] =8'h00;
         blockMem[173] =8'h00;
         blockMem[174] =8'h00;
         blockMem[175] =8'h00;
         blockMem[176] =8'h00;
         blockMem[177] =8'h00;
         blockMem[178] =8'h00;
         blockMem[179] =8'h00;
         blockMem[180] =8'h00;
         blockMem[181] =8'h00;
         blockMem[182] =8'h00;
         blockMem[183] =8'h00;
         blockMem[184] =8'h00;
         blockMem[185] =8'h00;
         blockMem[186] =8'h00;
         blockMem[187] =8'h00;
         blockMem[188] =8'h00;
         blockMem[189] =8'h00;
         blockMem[190] =8'h00;
         blockMem[191] =8'h00;
         blockMem[192] =8'h00;
         blockMem[193] =8'h00;
         blockMem[194] =8'h00;
         blockMem[195] =8'h00;
         blockMem[196] =8'h00;
         blockMem[197] =8'h00;
         blockMem[198] =8'h00;
         blockMem[199] =8'h00;
         blockMem[200] =8'h00;
         blockMem[201] =8'h00;
         blockMem[202] =8'h00;
         blockMem[203] =8'h00;
         blockMem[204] =8'h00;
         blockMem[205] =8'h00;
         blockMem[206] =8'h00;
         blockMem[207] =8'h00;
         blockMem[208] =8'h00;
         blockMem[209] =8'h00;
         blockMem[210] =8'h00;
         blockMem[211] =8'h00;
         blockMem[212] =8'h00;
         blockMem[213] =8'h00;
         blockMem[214] =8'h00;
         blockMem[215] =8'h00;
         blockMem[216] =8'h00;
         blockMem[217] =8'h00;
         blockMem[218] =8'h00;
         blockMem[219] =8'h00;
         blockMem[220] =8'h00;
         blockMem[221] =8'h00;
         blockMem[222] =8'h00;
         blockMem[223] =8'h00;
         blockMem[224] =8'h00;
         blockMem[225] =8'h00;
         blockMem[226] =8'h00;
         blockMem[227] =8'h00;
         blockMem[228] =8'h00;
         blockMem[229] =8'h00;
         blockMem[230] =8'h00;
         blockMem[231] =8'h00;
         blockMem[232] =8'h00;
         blockMem[233] =8'h00;
         blockMem[234] =8'h00;
         blockMem[235] =8'h00;
         blockMem[236] =8'h00;
         blockMem[237] =8'h00;
         blockMem[238] =8'h00;
         blockMem[239] =8'h00;
         blockMem[240] =8'h00;
         blockMem[241] =8'h00;
         blockMem[242] =8'h00;
         blockMem[243] =8'h00;
         blockMem[244] =8'h00;
         blockMem[245] =8'h00;
         blockMem[246] =8'h00;
         blockMem[247] =8'h00;
         blockMem[248] =8'h00;
         blockMem[249] =8'h00;
         blockMem[250] =8'h00;
         blockMem[251] =8'h00;
         blockMem[252] =8'h00;
         blockMem[253] =8'h00;
         blockMem[254] =8'h00;
         blockMem[255] =8'h00;     
    */
    end
endmodule
